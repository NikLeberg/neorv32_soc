-- =============================================================================
-- File:                    wb_imem.vhdl
--
-- Entity:                  wb_imem
--
-- Description:             Wishbone accessible instruction memory (IMEM).
--                          Implemented as dual-port ROM each port gets made
--                          accessible through one Wishbone slave channel. The
--                          idea is that two masters (i.e. CPUs) can access the
--                          instruction memory at the same time.
--
-- Note 1:                  Synthesizer should be inferring a synchronous dual-
--                          port ROM that gets used as RAM. Quartus Prime states
--                          successful inferring in a log message like so:
--                          "Info (19000): Inferred 1 megafunctions from design
--                          logic" and "Info (276031): Inferred altsyncram
--                          megafunction from the following design logic <>"
--
-- Note 2:                  Large chunks of this file are a 1:1 copy from
--                          neorv32_imem.default.vhd Copyright (c) 2023, Stephan
--                          Nolting. See respective file for more information.
--
-- Author:                  Niklaus Leuenberger <@NikLeberg>
--
-- SPDX-License-Identifier: MIT
--
-- Version:                 0.1
--
-- Changes:                 0.1, 2023-04-16, NikLeberg
--                              initial version
-- =============================================================================

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

LIBRARY neorv32;
USE neorv32.neorv32_package.ALL;
USE neorv32.neorv32_application_image.ALL; -- this file is generated by the image generator

USE work.wb_pkg.ALL;

ENTITY wb_imem IS
    GENERIC (
        IMEM_SIZE : NATURAL := 16 * 1024 -- size of instruction memory in bytes
    );
    PORT (
        -- Global control --
        clk_i  : IN STD_ULOGIC; -- global clock, rising edge
        rstn_i : IN STD_ULOGIC; -- global reset, low-active, sync

        -- Wishbone slave interfaces --
        wb_slaves_i : IN wb_req_arr_t(1 DOWNTO 0);  -- control and data from master to slave
        wb_slaves_o : OUT wb_resp_arr_t(1 DOWNTO 0) -- status and data from slave to master
    );
END ENTITY wb_imem;

ARCHITECTURE no_target_specific OF wb_imem IS

    -- application (image) size in bytes --
    CONSTANT imem_app_size_c : NATURAL := (application_init_image'length) * 4;

    -- ROM - initialized with executable code --
    CONSTANT mem_rom : mem32_t(0 TO IMEM_SIZE/4 - 1) := mem32_init_f(application_init_image, IMEM_SIZE/4);

    -- local signals --
    SIGNAL addr0, addr1 : STD_ULOGIC_VECTOR(index_size_f(IMEM_SIZE/4) - 1 DOWNTO 0);
    SIGNAL ack0, ack1, err0, err1 : STD_ULOGIC;

BEGIN

    -- Implement IMEM as pre-initialized dual-port ROM ----------------------------------------
    -- -------------------------------------------------------------------------------------------
    addr0 <= wb_slaves_i(0).adr(index_size_f(IMEM_SIZE/4) + 1 DOWNTO 2); -- word aligned
    addr1 <= wb_slaves_i(1).adr(index_size_f(IMEM_SIZE/4) + 1 DOWNTO 2); -- word aligned
    mem_access : PROCESS (clk_i)
    BEGIN
        IF rising_edge(clk_i) THEN
            -- Port A
            IF (wb_slaves_i(0).stb = '1') THEN -- reduce switching activity when not accessed
                wb_slaves_o(0).dat <= mem_rom(to_integer(unsigned(addr0)));
            END IF;
            -- Port B
            IF (wb_slaves_i(1).stb = '1') THEN -- reduce switching activity when not accessed
                wb_slaves_o(1).dat <= mem_rom(to_integer(unsigned(addr1)));
            END IF;
        END IF;
    END PROCESS mem_access;

    -- Bus Feedback ---------------------------------------------------------------------------
    -- -------------------------------------------------------------------------------------------
    bus_feedback : PROCESS (clk_i) IS
    BEGIN
        IF rising_edge(clk_i) THEN
            IF rstn_i = '0' THEN
                ack0 <= '0';
                err0 <= '0';
                ack1 <= '0';
                err1 <= '0';
            ELSE
                -- Ack' an access for one clock cycle only.
                IF wb_slaves_i(0).stb = '1' AND (ack0 OR err0) = '0' THEN
                    ack0 <= NOT wb_slaves_i(0).we;
                    err0 <= wb_slaves_i(0).we; -- read only!
                ELSE
                    ack0 <= '0';
                    err0 <= '0';
                END IF;
                IF wb_slaves_i(1).stb = '1' AND (ack1 OR err1) = '0' THEN
                    ack1 <= NOT wb_slaves_i(1).we;
                    err1 <= wb_slaves_i(1).we; -- read only!
                ELSE
                    ack1 <= '0';
                    err1 <= '0';
                END IF;
            END IF;
        END IF;
    END PROCESS bus_feedback;
    -- Master may abort the transmission, gate ack and err signals.
    wb_slaves_o(0).ack <= ack0 AND wb_slaves_i(0).stb;
    wb_slaves_o(0).err <= err0 AND wb_slaves_i(0).stb;
    wb_slaves_o(1).ack <= ack1 AND wb_slaves_i(1).stb;
    wb_slaves_o(1).err <= err1 AND wb_slaves_i(1).stb;

END ARCHITECTURE no_target_specific;
